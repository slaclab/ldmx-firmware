-------------------------------------------------------------------------------
-- Title      :
-------------------------------------------------------------------------------
-- Author     : Benjamin Reese  <bareese@slac.stanford.edu>
-------------------------------------------------------------------------------
-- Description:
-------------------------------------------------------------------------------
-- Copyright (c) 2013 SLAC National Accelerator Laboratory
-------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library UNISIM;
use UNISIM.VCOMPONENTS.all;


library surf;
use surf.StdRtlPkg.all;
use surf.AxiLitePkg.all;
use surf.AxiStreamPkg.all;
use surf.Pgp2FcPkg.all;

library lcls_timing_core;
use lcls_timing_core.TimingPkg.all;

library ldmx_tdaq;
use ldmx_tdaq.FcPkg.all;

entity FcHub is

   generic (
      TPD_G             : time                 := 1 ns;
      SIM_SPEEDUP_G     : boolean              := false;
      REFCLKS_G         : integer range 1 to 4 := 1;
      QUADS_G           : integer range 1 to 4 := 1;
      QUAD_REFCLK_MAP_G : IntegerArray         := (0      => 0);  --, 1 => 0, 2 => 1, 3 => 1);  -- Map a refclk for each quad
      AXIL_CLK_FREQ_G   : real                 := 156.25e6;
      AXIL_BASE_ADDR_G  : slv(31 downto 0)     := (others => '0'));
   port (
      ----------------------------------------------------------------------------------------------
      -- LCLS Timing Interface
      ----------------------------------------------------------------------------------------------
      -- 185/371 MHz Ref Clk for LCLS timing recovery (freq used depends on GT configuration)
      lclsTimingRefClkP : in  sl;
      lclsTimingRefClkN : in  sl;
      -- LCLS-II timing interface
      lclsTimingRxP     : in  sl;
      lclsTimingRxN     : in  sl;
      lclsTimingTxP     : out sl;
      lclsTimingTxN     : out sl;
      -- Recovered clock via GT dedicated clock pins
      timingRecClkOutP  : out sl;
      timingRecClkOutN  : out sl;

      ----------------------------------------------------------------------------------------------
      -- Global Trigger Interface
      ----------------------------------------------------------------------------------------------
      -- LCLS Recovered Clock Output via fabric pins
      lclsTimingClkOut  : out sl;
      lclsTimingRstOut  : out sl;
      lclsTimingFcTxMsg : out FcMessageType;
      lclsTimingBus     : out TimingBusType;
      globalTriggerRor  : in  FcTimestampType;

      ----------------------------------------------------------------------------------------------
      -- FC HUB
      ----------------------------------------------------------------------------------------------
      -- Recovered and retimed LCLS Reference clock
      fcHubRefClkP : in  slv(REFCLKS_G-1 downto 0);
      fcHubRefClkN : in  slv(REFCLKS_G-1 downto 0);
      -- PGP FC serial IO
      fcHubTxP     : out slv(QUADS_G*4-1 downto 0);
      fcHubTxN     : out slv(QUADS_G*4-1 downto 0);
      fcHubRxP     : in  slv(QUADS_G*4-1 downto 0);
      fcHubRxN     : in  slv(QUADS_G*4-1 downto 0);

      ----------------------------------------------------------------------------------------------
      -- AXI Lite
      ----------------------------------------------------------------------------------------------
      axilClk         : in  sl;
      axilRst         : in  sl;
      axilReadMaster  : in  AxiLiteReadMasterType;
      axilReadSlave   : out AxiLiteReadSlaveType;
      axilWriteMaster : in  AxiLiteWriteMasterType;
      axilWriteSlave  : out AxiLiteWriteSlaveType);

end entity FcHub;

architecture rtl of FcHub is

   -- AXI Lite
   constant AXIL_NUM_C         : integer := 3;
   constant AXIL_LCLS_TIMING_C : integer := 0;
   constant AXIL_TX_LOGIC_C    : integer := 1;
   constant AXIL_FC_ARRAY_C    : integer := 2;

   constant AXIL_XBAR_CONFIG_C : AxiLiteCrossbarMasterConfigArray(AXIL_NUM_C-1 downto 0) := (
      AXIL_LCLS_TIMING_C => (
         baseAddr        => AXIL_BASE_ADDR_G + X"0000_0000",
         addrBits        => 20,
         connectivity    => X"FFFF"),
      AXIL_TX_LOGIC_C    => (
         baseAddr        => AXIL_BASE_ADDR_G +X"0010_0000",
         addrBits        => 8,
         connectivity    => X"FFFF"),
      AXIL_FC_ARRAY_C    => (
         baseAddr        => AXIL_BASE_ADDR_G +X"0020_0000",
         addrBits        => 20,
         connectivity    => X"FFFF"));

   signal locAxilReadMasters  : AxiLiteReadMasterArray(AXIL_NUM_C-1 downto 0);
   signal locAxilReadSlaves   : AxiLiteReadSlaveArray(AXIL_NUM_C-1 downto 0)  := (others => AXI_LITE_READ_SLAVE_EMPTY_DECERR_C);
   signal locAxilWriteMasters : AxiLiteWriteMasterArray(AXIL_NUM_C-1 downto 0);
   signal locAxilWriteSlaves  : AxiLiteWriteSlaveArray(AXIL_NUM_C-1 downto 0) := (others => AXI_LITE_WRITE_SLAVE_EMPTY_DECERR_C);

   -- Recovered LCLS Timing Clock and Bus
   signal lclsTimingClk    : sl;
   signal lclsTimingRst    : sl;
   signal lclsTimingBusLoc : TimingBusType;

   -- LDMX Fast Control Message to FC Senders
   signal fcTxMsg : FcMessageType;

begin

   -------------------------------------------------------------------------------------------------
   -- AXI-Lite crossbar
   -------------------------------------------------------------------------------------------------
   U_XBAR : entity surf.AxiLiteCrossbar
      generic map (
         TPD_G              => TPD_G,
         NUM_SLAVE_SLOTS_G  => 1,
         NUM_MASTER_SLOTS_G => AXIL_NUM_C,
         MASTERS_CONFIG_G   => AXIL_XBAR_CONFIG_C)
      port map (
         axiClk              => axilClk,
         axiClkRst           => axilRst,
         sAxiWriteMasters(0) => axilWriteMaster,
         sAxiWriteSlaves(0)  => axilWriteSlave,
         sAxiReadMasters(0)  => axilReadMaster,
         sAxiReadSlaves(0)   => axilReadSlave,
         mAxiWriteMasters    => locAxilWriteMasters,
         mAxiWriteSlaves     => locAxilWriteSlaves,
         mAxiReadMasters     => locAxilReadMasters,
         mAxiReadSlaves      => locAxilReadSlaves);


   -------------------------------------------------------------------------------------------------
   -- LCLS TIMING RX
   -------------------------------------------------------------------------------------------------
   lclsTimingClkOut <= lclsTimingClk;
   lclsTimingBus    <= lclsTimingBusLoc;

   U_Lcls2TimingRx_1 : entity ldmx_tdaq.Lcls2TimingRx
      generic map (
         TPD_G             => TPD_G,
         SIMULATION_G      => SIM_SPEEDUP_G,
         TIME_GEN_EXTREF_G => true,
         RX_CLK_MMCM_G     => true,
         USE_TPGMINI_G     => true,
         AXI_CLK_FREQ_G    => AXIL_CLK_FREQ_G,
         AXIL_BASE_ADDR_G  => AXIL_XBAR_CONFIG_C(AXIL_LCLS_TIMING_C).baseAddr)
      port map (
         stableClk        => axilClk,   -- [in] -- axilClk from TenGigEth core is not mmcm
         stableRst        => axilRst,   -- [in]
         axilClk          => axilClk,   -- [in]
         axilRst          => axilRst,   -- [in]
         axilReadMaster   => locAxilReadMasters(AXIL_LCLS_TIMING_C),   -- [in]
         axilReadSlave    => locAxilReadSlaves(AXIL_LCLS_TIMING_C),    -- [out]
         axilWriteMaster  => locAxilWriteMasters(AXIL_LCLS_TIMING_C),  -- [in]
         axilWriteSlave   => locAxilWriteSlaves(AXIL_LCLS_TIMING_C),   -- [out]
         recTimingClk     => lclsTimingClk,                            -- [out]
         recTimingRst     => lclsTimingRst,                            -- [out]
         appTimingBus     => lclsTimingBusLoc,                         -- [out]
         timingRxP        => lclsTimingRxP,                            -- [in]
         timingRxN        => lclsTimingRxN,                            -- [in]
         timingTxP        => lclsTimingTxP,                            -- [out]
         timingTxN        => lclsTimingTxN,                            -- [out]
         timingRefClkInP  => lclsTimingRefClkP,                        -- [in]
         timingRefClkInN  => lclsTimingRefClkN,                        -- [in]
         timingRecClkOutP => timingRecClkOutP,                         -- [out]
         timingRecClkOutN => timingRecClkOutN);                        -- [out]

   -------------------------------------------------------------------------------------------------
   -- Fast Control Output Word Logic
   -------------------------------------------------------------------------------------------------
   U_FcTxLogic_1 : entity ldmx_tdaq.FcTxLogic
      generic map (
         TPD_G => TPD_G)
      port map (
         lclsTimingClk    => lclsTimingClk,                         -- [in]
         lclsTimingRst    => lclsTimingRst,                         -- [in]
         lclsTimingBus    => lclsTimingBusLoc,                      -- [in]
         globalTriggerRor => globalTriggerRor,                      -- [in]
         fcMsg            => fcTxMsg,                               -- [out]
         axilClk          => axilClk,                               -- [in]
         axilRst          => axilRst,                               -- [in]
         axilReadMaster   => locAxilReadMasters(AXIL_TX_LOGIC_C),   -- [in]
         axilReadSlave    => locAxilReadSlaves(AXIL_TX_LOGIC_C),    -- [out]
         axilWriteMaster  => locAxilWriteMasters(AXIL_TX_LOGIC_C),  -- [in]
         axilWriteSlave   => locAxilWriteSlaves(AXIL_TX_LOGIC_C));  -- [out]

   -------------------------------------------------------------------------------------------------
   -- Fast Control Fanout to Subsystems
   -------------------------------------------------------------------------------------------------
   U_FcSenderArray_1 : entity ldmx_tdaq.FcSenderArray
      generic map (
         TPD_G             => TPD_G,
         SIM_SPEEDUP_G     => SIM_SPEEDUP_G,
         REFCLKS_G         => REFCLKS_G,
         QUADS_G           => QUADS_G,
         QUAD_REFCLK_MAP_G => QUAD_REFCLK_MAP_G,
         AXIL_CLK_FREQ_G   => AXIL_CLK_FREQ_G,
         AXIL_BASE_ADDR_G  => AXIL_XBAR_CONFIG_C(AXIL_FC_ARRAY_C).baseAddr)
      port map (
         fcHubRefClkP    => fcHubRefClkP,                          -- [in]
         fcHubRefClkN    => fcHubRefClkN,                          -- [in]
         fcHubTxP        => fcHubTxP,                              -- [out]
         fcHubTxN        => fcHubTxN,                              -- [out]
         fcHubRxP        => fcHubRxP,                              -- [in]
         fcHubRxN        => fcHubRxN,                              -- [in]
         lclsTimingClk   => lclsTimingClk,                         -- [in]
         lclsTimingRst   => lclsTimingRst,                         -- [in]
         fcTxMsg         => fcTxMsg,                               -- [in]
         axilClk         => axilClk,                               -- [in]
         axilRst         => axilRst,                               -- [in]
         axilReadMaster  => locAxilReadMasters(AXIL_FC_ARRAY_C),   -- [in]
         axilReadSlave   => locAxilReadSlaves(AXIL_FC_ARRAY_C),    -- [out]
         axilWriteMaster => locAxilWriteMasters(AXIL_FC_ARRAY_C),  -- [in]
         axilWriteSlave  => locAxilWriteSlaves(AXIL_FC_ARRAY_C));  -- [out]


end rtl;
